module top_module( 
    input a, 
    input b, 
    output out );
    
    reg out1;
    
    assign out1 = a^b;
    assign out = ~out1;

endmodule
